module cpu_top (
    input clk,
    input reset_n


);

wire redirect_valid;
wire [31:0] redirect_target_pc;

endmodule